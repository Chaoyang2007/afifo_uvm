`include "uvm_macros.svh"

import uvm_pkg::*;
